library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity subBytes is
    port (
	 clock    : std_logic;
    address  : in std_logic_Vector(7 downto 0);
    data     : out std_logic_Vector(7 downto 0)
    );
end subBytes;

architecture  rtl of subBytes is

  type mem is array (0 to 255) of std_logic_vector(7 downto 0);
     constant my_Rom : mem := (
			0  => "01100011",
			1  => "01111100",
			2  => "01110111",
			3  => "01111011",
			4  => "11110010",
			5  => "01101011",
			6  => "01101111",
			7  => "11000101",
			8  => "11000101",
			9  => "00000001",
			10 => "01100111",
			11 => "00101011",
			12 => "11111110",
			13 => "11010111",
			14 => "10101011",
			15 => "01110110",
			16 => "11001010",
			17 => "10000010",
			18 => "11001001",
			19 => "01111101",
			20 => "11111010",
			21 => "01011001",
			22 => "01000111",
			23 => "11110000",
			24 => "10101101",
			25 => "11010100",
			26 => "10100010",
			27 => "10101111",
			28 => "10011100",
			29 => "10100100",
			30 => "01110010",
			31 => "11000000",
			32 => "10110111",
			33 => "11111101",
			34 => "10010011",
			35 => "00100110",
			36 => "00110110",
			37 => "00111111",
			38 => "11110111",
			39 => "11001100",
			40 => "00110100",
			41 => "10100101",
			42 => "11100101", 
			43 => "11110001",
			44 => "01110001",
			45 => "11011000", 
			46 => "00110001",
			47 => "00010101",
			48 => "00000100",
			49 => "11000111",
			50 => "00100011",
			51 => "11000011",
			52 => "00011000",
			53 => "10010110",
			54 => "00000101",
			55 => "10011010",
			56 => "00000111",
			57 => "00010010",
			58 => "10000000",
			59 => "11100010",
			60 => "11101011",
			61 => "00100111",
			62 => "10110010",
			63 => "01110101",
			64 => "00001001",
			65 => "10000011",
			66 => "00101100",
			67 => "00011010",
			68 => "00011011", 
			69 => "01101110",
			70 => "01011010",
			71 => "10100000",
			72 => "01010010",
			73 => "00111011",
			74 => "11010110",
			75 => "10110011",
			76 => "00101001",
			77 => "11100011",
			78 => "00101111",
			79 => "10000100",
			80 => "01010011",
			81 => "11010001",
			82 => "00000000",
			83 => "11101101",
			84 => "00100000",
			85 => "11111100",
			86 => "10110001", 
			87 => "01011011", 
			88 => "01101010",
			89 => "11001011", 
			90 => "10111110",
			91 => "00111001",
			92 => "01001010",
			93 => "01001100",
			94 => "01011000", 
			95 => "11001111",
			96 => "11010000", 
			97 => "11101111",
			98 => "10101010",
			99 => "11111011",
			100 => "01000011",
			101 => "01001101",
			102 => "00110011", 
			103 => "10000101",
			104 => "01000101",
			105 => "11111001",
			106 => "00000010", 
			107 => "01111111",
			108 => "01010000",
			109 => "00111100",
			110 => "00111100",
			111 => "10101000",
			112 => "01010001",
			113 => "10100011",
			114 => "01000000",
			115 => "10001111",
			116 => "10010010",
			117 => "10011101",
			118 => "00111000",
			119 => "11110101",
			120 => "10111100", 
			121 => "10110110",
			122 => "11011010",
			123 => "00100001",
			124 => "00010000",
			125 => "11111111",
			126 => "11110011",
			127 => "11010010",
			128 => "11001101",
			129 => "00001100",
			130 => "00010011",
			131 => "11101100",
			132 => "01011111",
			133 => "10010111",
			134 => "01000100",
			135 => "00010111",
			136 => "11000100",
			137 => "10100111",
			138 => "01111110",
			139 => "00111101",
			140 => "01100100",
			141 => "01100100",
			142 => "00011001",
			143 => "01110011",
			144 => "01100000",
			145 => "10000001",
			146 => "01001111",
			147 => "11011100", 
			148 => "00100010",
			149 => "00101010",
			150 => "10010000",
			151 => "10001000",
			152 => "01000110",
			153 => "11101110",
			154 => "10111000",
			155 => "00010100",
			156 => "11011110",
			157 => "01011110",
			158 => "00001011",
			159 => "11011011",
			160 => "11100000",
			161 => "00110010",
			162 => "00111010",
			163 => "00001010",
			164 => "01001001", 
			165 => "00000110",
			166 => "00100100",
			167 => "01011100",
			168 => "11000010",
			169 => "11010011",
			170 => "10101100",
			171 => "01100010",
			172 => "10010001",
			173 => "10010101",
			174 => "11100100",
			175 => "01111001",
			176 => "11100111",
			177 => "11001000",
			178 => "00110111",
			179 => "01101101",
			180 => "10001101",
			181 => "11010101",
			182 => "01001110",
			183 => "10101001",
			184 => "01101100",
			185 => "01010110", 
			186 => "11110100",
			187 => "11101010", 
			188 => "01100101",
			189 => "01111010",
			190 => "10101110",
			191 => "00001000",
			192 => "10111010",
			193 => "01111000",
			194 => "00100101",
			195 => "00101110",
			196 => "00011100",
			197 => "10100110",
			198 => "10110100",
			199 => "11000110",
			200 => "11101000",
			201 => "11011101",
			202 => "01110100", 
			203 => "00001111",
			204 => "01001011",
			205 => "10111101",
			206 => "10001011",
			207 => "10001010",
			208 => "01110000", 
			209 => "00111110",
			210 => "10110101", 
			211 => "01100110",
			212 => "01001000",
			213 => "00000011",
			214 => "11110110",
			215 => "00001110",
			216 => "01100001",
			217 => "00110101",
			218 => "01010111",
			219 => "10111001",
			220 => "10000110",
			221 => "11000001",
			222 => "00011101", 
			223 => "10011110",
			224 => "11100001",
			225 => "11111000",
			226 => "10011000",
			227 => "00010001",
			228 => "01101001", 
			229 => "11011001",
			230 => "10001110",
			231 => "10010100", 
			232 => "10011011",
			233 => "00011110",
			234 => "10000111",
			235 => "11101001",
			236 => "11001110",
			237 => "01010101",
			238 => "00101000",
			239 => "11011111",
			240 => "10001100",
			241 => "10100001",
			242 => "10001001",
			243 => "00001101",
			244 => "10111111",
			245 => "11100110",
			246 => "01000010",
			247 => "01101000", 
			248 => "01000001",
			249 => "10011001",
			250 => "00101101",
			251 => "00001111",
			252 => "10110000",
			253 => "01010100",
			254 => "01010100",
			255 => "00010110"
       );



begin
  process (address)
  begin
    case address is
      when "00000000" => data <= my_rom(0);
		when "00000001" => data <= my_rom(1);
		when "00000010" => data <= my_rom(2);
		when "00000011" => data <= my_rom(3);
		when "00000100" => data <= my_rom(4);
		when "00000101" => data <= my_rom(5);
		when "00000110" => data <= my_rom(6);
		when "00000111" => data <= my_rom(7);
		when "00001000" => data <= my_rom(8);
		when "00001001" => data <= my_rom(9);
		when "00001010" => data <= my_rom(10);
		when "00001011" => data <= my_rom(11);
		when "00001100" => data <= my_rom(12);
		when "00001101" => data <= my_rom(13);
		when "00001110" => data <= my_rom(14);
		when "00001111" => data <= my_rom(15);
		when "00010000" => data <= my_rom(16);
		when "00010001" => data <= my_rom(17);
		when "00010010" => data <= my_rom(18);
		when "00010011" => data <= my_rom(19);
		when "00010100" => data <= my_rom(20);
		when "00010101" => data <= my_rom(21);
		when "00010110" => data <= my_rom(22);
		when "00010111" => data <= my_rom(23);
		when "00011000" => data <= my_rom(24);
		when "00011001" => data <= my_rom(25);
		when "00011010" => data <= my_rom(26);
		when "00011011" => data <= my_rom(27);
		when "00011100" => data <= my_rom(28);
		when "00011101" => data <= my_rom(29);
		when "00011110" => data <= my_rom(30);
		when "00011111" => data <= my_rom(31);
		when "00100000" => data <= my_rom(32);
		when "00100001" => data <= my_rom(33);
		when "00100010" => data <= my_rom(34);
		when "00100011" => data <= my_rom(35);
		when "00100100" => data <= my_rom(36);
		when "00100101" => data <= my_rom(37);
		when "00100110" => data <= my_rom(38);
		when "00100111" => data <= my_rom(39);
		when "00101000" => data <= my_rom(40);
		when "00101001" => data <= my_rom(41);
		when "00101010" => data <= my_rom(42);
		when "00101011" => data <= my_rom(43);
		when "00101100" => data <= my_rom(44);
		when "00101101" => data <= my_rom(45);
		when "00101110" => data <= my_rom(46);
		when "00101111" => data <= my_rom(47);
		when "00110000" => data <= my_rom(48);
		when "00110001" => data <= my_rom(49);
		when "00110010" => data <= my_rom(50);
		when "00110011" => data <= my_rom(51);
		when "00110100" => data <= my_rom(52);
		when "00110101" => data <= my_rom(53);
		when "00110110" => data <= my_rom(54);
		when "00110111" => data <= my_rom(55);
		when "00111000" => data <= my_rom(56);
		when "00111001" => data <= my_rom(57);
		when "00111010" => data <= my_rom(58);
		when "00111011" => data <= my_rom(59);
		when "00111100" => data <= my_rom(60);
		when "00111101" => data <= my_rom(61);
		when "00111110" => data <= my_rom(62);
		when "00111111" => data <= my_rom(63);
		when "01000000" => data <= my_rom(64);
		when "01000001" => data <= my_rom(65);
		when "01000010" => data <= my_rom(66);
		when "01000011" => data <= my_rom(67);
		when "01000100" => data <= my_rom(68);
		when "01000101" => data <= my_rom(69);
		when "01000110" => data <= my_rom(70);
		when "01000111" => data <= my_rom(71);
		when "01001000" => data <= my_rom(72);
		when "01001001" => data <= my_rom(73);
		when "01001010" => data <= my_rom(74);
		when "01001011" => data <= my_rom(75);
		when "01001100" => data <= my_rom(76);
		when "01001101" => data <= my_rom(77);
		when "01001110" => data <= my_rom(78);
		when "01001111" => data <= my_rom(79);
		when "01010000" => data <= my_rom(80);
		when "01010001" => data <= my_rom(81);
		when "01010010" => data <= my_rom(82);
		when "01010011" => data <= my_rom(83);
		when "01010100" => data <= my_rom(84);
		when "01010101" => data <= my_rom(85);
		when "01010110" => data <= my_rom(86);
		when "01010111" => data <= my_rom(87);
		when "01011000" => data <= my_rom(88);
		when "01011001" => data <= my_rom(89);
		when "01011010" => data <= my_rom(90);
		when "01011011" => data <= my_rom(91);
		when "01011100" => data <= my_rom(92);
		when "01011101" => data <= my_rom(93);
		when "01011110" => data <= my_rom(94);
		when "01011111" => data <= my_rom(95);
		when "01100000" => data <= my_rom(96);
		when "01100001" => data <= my_rom(97);
		when "01100010" => data <= my_rom(98);
		when "01100011" => data <= my_rom(99);
		when "01100100" => data <= my_rom(100);
		when "01100101" => data <= my_rom(101);
		when "01100110" => data <= my_rom(102);
		when "01100111" => data <= my_rom(103);
		when "01101000" => data <= my_rom(104);
		when "01101001" => data <= my_rom(105);
		when "01101010" => data <= my_rom(106);
		when "01101011" => data <= my_rom(107);
		when "01101100" => data <= my_rom(108);
		when "01101101" => data <= my_rom(109);
		when "01101110" => data <= my_rom(110);
		when "01101111" => data <= my_rom(111);
		when "01110000" => data <= my_rom(112);
		when "01110001" => data <= my_rom(113);
		when "01110010" => data <= my_rom(114);
		when "01110011" => data <= my_rom(115);
		when "01110100" => data <= my_rom(116);
		when "01110101" => data <= my_rom(117);
		when "01110110" => data <= my_rom(118);
		when "01110111" => data <= my_rom(119);
		when "01111000" => data <= my_rom(120);
		when "01111001" => data <= my_rom(121);
		when "01111010" => data <= my_rom(122);
		when "01111011" => data <= my_rom(123);
		when "01111100" => data <= my_rom(124);
		when "01111101" => data <= my_rom(125);
		when "01111110" => data <= my_rom(126);
		when "01111111" => data <= my_rom(127);
		when "10000000" => data <= my_rom(128);
		when "10000001" => data <= my_rom(129);
		when "10000010" => data <= my_rom(130);
		when "10000011" => data <= my_rom(131);
		when "10000100" => data <= my_rom(132);
		when "10000101" => data <= my_rom(133);
		when "10000110" => data <= my_rom(134);
		when "10000111" => data <= my_rom(135);
		when "10001000" => data <= my_rom(136);
		when "10001001" => data <= my_rom(137);
		when "10001010" => data <= my_rom(138);
		when "10001011" => data <= my_rom(139);
		when "10001100" => data <= my_rom(140);
		when "10001101" => data <= my_rom(141);
		when "10001110" => data <= my_rom(142);
		when "10001111" => data <= my_rom(143);
		when "10010000" => data <= my_rom(144);
		when "10010001" => data <= my_rom(145);
		when "10010010" => data <= my_rom(146);
		when "10010011" => data <= my_rom(147);
		when "10010100" => data <= my_rom(148);
		when "10010101" => data <= my_rom(149);
		when "10010110" => data <= my_rom(150);
		when "10010111" => data <= my_rom(151);
		when "10011000" => data <= my_rom(152);
		when "10011001" => data <= my_rom(153);
		when "10011010" => data <= my_rom(154);
		when "10011011" => data <= my_rom(155);
		when "10011100" => data <= my_rom(156);
		when "10011101" => data <= my_rom(157);
		when "10011110" => data <= my_rom(158);
		when "10011111" => data <= my_rom(159);
		when "10100000" => data <= my_rom(160);
		when "10100001" => data <= my_rom(161);
		when "10100010" => data <= my_rom(162);
		when "10100011" => data <= my_rom(163);
		when "10100100" => data <= my_rom(164);
		when "10100101" => data <= my_rom(165);
		when "10100110" => data <= my_rom(166);
		when "10100111" => data <= my_rom(167);
		when "10101000" => data <= my_rom(168);
		when "10101001" => data <= my_rom(169);
		when "10101010" => data <= my_rom(170);
		when "10101011" => data <= my_rom(171);
		when "10101100" => data <= my_rom(172);
		when "10101101" => data <= my_rom(173);
		when "10101110" => data <= my_rom(174);
		when "10101111" => data <= my_rom(175);
		when "10110000" => data <= my_rom(176);
		when "10110001" => data <= my_rom(177);
		when "10110010" => data <= my_rom(178);
		when "10110011" => data <= my_rom(179);
		when "10110100" => data <= my_rom(180);
		when "10110101" => data <= my_rom(181);
		when "10110110" => data <= my_rom(182);
		when "10110111" => data <= my_rom(183);
		when "10111000" => data <= my_rom(184);
		when "10111001" => data <= my_rom(185);
		when "10111010" => data <= my_rom(186);
		when "10111011" => data <= my_rom(187);
		when "10111100" => data <= my_rom(188);
		when "10111101" => data <= my_rom(189);
		when "10111110" => data <= my_rom(190);
		when "10111111" => data <= my_rom(191);
		when "11000000" => data <= my_rom(192);
		when "11000001" => data <= my_rom(193);
		when "11000010" => data <= my_rom(194);
		when "11000011" => data <= my_rom(195);
		when "11000100" => data <= my_rom(196);
		when "11000101" => data <= my_rom(197);
		when "11000110" => data <= my_rom(198);
		when "11000111" => data <= my_rom(199);
		when "11001000" => data <= my_rom(200);
		when "11001001" => data <= my_rom(201);
		when "11001010" => data <= my_rom(202);
		when "11001011" => data <= my_rom(203);
		when "11001100" => data <= my_rom(204);
		when "11001101" => data <= my_rom(205);
		when "11001110" => data <= my_rom(206);
		when "11001111" => data <= my_rom(207);
		when "11010000" => data <= my_rom(208);
		when "11010001" => data <= my_rom(209);
		when "11010010" => data <= my_rom(210);
		when "11010011" => data <= my_rom(211);
		when "11010100" => data <= my_rom(212);
		when "11010101" => data <= my_rom(213);
		when "11010110" => data <= my_rom(214);
		when "11010111" => data <= my_rom(215);
		when "11011000" => data <= my_rom(216);
		when "11011001" => data <= my_rom(217);
		when "11011010" => data <= my_rom(218);
		when "11011011" => data <= my_rom(219);
		when "11011100" => data <= my_rom(220);
		when "11011101" => data <= my_rom(221);
		when "11011110" => data <= my_rom(222);
		when "11011111" => data <= my_rom(223);
		when "11100000" => data <= my_rom(224);
		when "11100001" => data <= my_rom(225);
		when "11100010" => data <= my_rom(226);
		when "11100011" => data <= my_rom(227);
		when "11100100" => data <= my_rom(228);
		when "11100101" => data <= my_rom(229);
		when "11100110" => data <= my_rom(230);
		when "11100111" => data <= my_rom(231);
		when "11101000" => data <= my_rom(232);
		when "11101001" => data <= my_rom(233);
		when "11101010" => data <= my_rom(234);
		when "11101011" => data <= my_rom(235);
		when "11101100" => data <= my_rom(236);
		when "11101101" => data <= my_rom(237);
		when "11101110" => data <= my_rom(238);
		when "11101111" => data <= my_rom(239);
		when "11110000" => data <= my_rom(240);
		when "11110001" => data <= my_rom(241);
		when "11110010" => data <= my_rom(242);
		when "11110011" => data <= my_rom(243);
		when "11110100" => data <= my_rom(244);
		when "11110101" => data <= my_rom(245);
		when "11110110" => data <= my_rom(246);
		when "11110111" => data <= my_rom(247);
		when "11111000" => data <= my_rom(248);
		when "11111001" => data <= my_rom(249);
		when "11111010" => data <= my_rom(250);
		when "11111011" => data <= my_rom(251);
		when "11111100" => data <= my_rom(252);
		when "11111101" => data <= my_rom(253);
		when "11111110" => data <= my_rom(254);
		when "11111111" => data <= my_rom(255);
  end case;
 end process;

end architecture;